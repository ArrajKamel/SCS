library ieee; 
use ieee.std_logic_1164.all; 
use ieee.unsigned_arith.all; 

entity carry_lookahead_adder is 
    port(
        
    );